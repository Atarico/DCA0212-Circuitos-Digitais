library verilog;
use verilog.vl_types.all;
entity mux4_in4bits_vlg_check_tst is
    port(
        saidam          : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end mux4_in4bits_vlg_check_tst;
