library verilog;
use verilog.vl_types.all;
entity hex7segdecode_vlg_vec_tst is
end hex7segdecode_vlg_vec_tst;
