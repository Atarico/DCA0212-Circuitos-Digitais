library verilog;
use verilog.vl_types.all;
entity display7seg_vlg_vec_tst is
end display7seg_vlg_vec_tst;
