library verilog;
use verilog.vl_types.all;
entity mux4_in4bits_vlg_vec_tst is
end mux4_in4bits_vlg_vec_tst;
